magic
tech sky130A
magscale 1 2
timestamp 1636924791
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 14 2128 199902 197520
<< metal2 >>
rect 32218 199200 32274 200000
rect 88154 199200 88210 200000
rect 144090 199200 144146 200000
rect 199842 199200 199898 200000
rect 18 0 74 800
rect 55770 0 55826 800
rect 111706 0 111762 800
rect 167642 0 167698 800
<< obsm2 >>
rect 20 199144 32162 199200
rect 32330 199144 88098 199200
rect 88266 199144 144034 199200
rect 144202 199144 199786 199200
rect 20 856 199896 199144
rect 130 800 55714 856
rect 55882 800 111650 856
rect 111818 800 167586 856
rect 167754 800 199896 856
<< metal3 >>
rect 0 165112 800 165232
rect 199200 117240 200000 117360
rect 0 82424 800 82544
rect 199200 34552 200000 34672
<< obsm3 >>
rect 800 165312 199200 197505
rect 880 165032 199200 165312
rect 800 117440 199200 165032
rect 800 117160 199120 117440
rect 800 82624 199200 117160
rect 880 82344 199200 82624
rect 800 34752 199200 82344
rect 800 34472 199120 34752
rect 800 2143 199200 34472
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< labels >>
rlabel metal3 s 0 82424 800 82544 6 CLK
port 1 nsew signal input
rlabel metal2 s 199842 199200 199898 200000 6 OUT[0]
port 2 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 OUT[1]
port 3 nsew signal output
rlabel metal2 s 18 0 74 800 6 OUT[2]
port 4 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 OUT[3]
port 5 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 OUT[4]
port 6 nsew signal output
rlabel metal2 s 144090 199200 144146 200000 6 OUT[5]
port 7 nsew signal output
rlabel metal3 s 199200 117240 200000 117360 6 OUT[6]
port 8 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 OUT[7]
port 9 nsew signal output
rlabel metal2 s 32218 199200 32274 200000 6 OUT[8]
port 10 nsew signal output
rlabel metal2 s 88154 199200 88210 200000 6 OUT[9]
port 11 nsew signal output
rlabel metal3 s 199200 34552 200000 34672 6 reset
port 12 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 13 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 14 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 14 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 14 nsew ground input
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 14 nsew ground input
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 14 nsew ground input
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 14 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 31821524
string GDS_START 761774
<< end >>

