magic
tech sky130A
magscale 1 2
timestamp 1636718384
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 14 2128 299998 297616
<< metal2 >>
rect 48410 299200 48466 300000
rect 132314 299200 132370 300000
rect 216218 299200 216274 300000
rect 299938 299200 299994 300000
rect 18 0 74 800
rect 83738 0 83794 800
rect 167642 0 167698 800
rect 251546 0 251602 800
<< obsm2 >>
rect 20 299144 48354 299200
rect 48522 299144 132258 299200
rect 132426 299144 216162 299200
rect 216330 299144 299882 299200
rect 20 856 299992 299144
rect 130 800 83682 856
rect 83850 800 167586 856
rect 167754 800 251490 856
rect 251658 800 299992 856
<< metal3 >>
rect 0 247800 800 247920
rect 299200 175992 300000 176112
rect 0 123768 800 123888
rect 299200 51960 300000 52080
<< obsm3 >>
rect 800 248000 299200 297601
rect 880 247720 299200 248000
rect 800 176192 299200 247720
rect 800 175912 299120 176192
rect 800 123968 299200 175912
rect 880 123688 299200 123968
rect 800 52160 299200 123688
rect 800 51880 299120 52160
rect 800 2143 299200 51880
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 142848 115635 157728 211309
rect 158208 115635 173088 211309
rect 173568 115635 183941 211309
<< labels >>
rlabel metal3 s 0 123768 800 123888 6 CLK
port 1 nsew signal input
rlabel metal2 s 299938 299200 299994 300000 6 OUT[0]
port 2 nsew signal output
rlabel metal3 s 0 247800 800 247920 6 OUT[1]
port 3 nsew signal output
rlabel metal2 s 18 0 74 800 6 OUT[2]
port 4 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 OUT[3]
port 5 nsew signal output
rlabel metal2 s 251546 0 251602 800 6 OUT[4]
port 6 nsew signal output
rlabel metal2 s 216218 299200 216274 300000 6 OUT[5]
port 7 nsew signal output
rlabel metal3 s 299200 175992 300000 176112 6 OUT[6]
port 8 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 OUT[7]
port 9 nsew signal output
rlabel metal2 s 48410 299200 48466 300000 6 OUT[8]
port 10 nsew signal output
rlabel metal2 s 132314 299200 132370 300000 6 OUT[9]
port 11 nsew signal output
rlabel metal3 s 299200 51960 300000 52080 6 reset
port 12 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 13 nsew power input
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 14 nsew ground input
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 14 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 300000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 44914778
string GDS_START 742720
<< end >>

