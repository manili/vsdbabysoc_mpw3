VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END CLK
  PIN OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 1496.000 1499.970 1500.000 ;
    END
  END OUT[0]
  PIN OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.000 4.000 1239.600 ;
    END
  END OUT[1]
  PIN OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END OUT[2]
  PIN OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END OUT[3]
  PIN OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.730 0.000 1258.010 4.000 ;
    END
  END OUT[4]
  PIN OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 1496.000 1081.370 1500.000 ;
    END
  END OUT[5]
  PIN OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 879.960 1500.000 880.560 ;
    END
  END OUT[6]
  PIN OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END OUT[7]
  PIN OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 1496.000 242.330 1500.000 ;
    END
  END OUT[8]
  PIN OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 1496.000 661.850 1500.000 ;
    END
  END OUT[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 259.800 1500.000 260.400 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 1499.990 1488.080 ;
      LAYER met2 ;
        RECT 0.100 1495.720 241.770 1496.000 ;
        RECT 242.610 1495.720 661.290 1496.000 ;
        RECT 662.130 1495.720 1080.810 1496.000 ;
        RECT 1081.650 1495.720 1499.410 1496.000 ;
        RECT 0.100 4.280 1499.960 1495.720 ;
        RECT 0.650 4.000 418.410 4.280 ;
        RECT 419.250 4.000 837.930 4.280 ;
        RECT 838.770 4.000 1257.450 4.280 ;
        RECT 1258.290 4.000 1499.960 4.280 ;
      LAYER met3 ;
        RECT 4.000 1240.000 1496.000 1488.005 ;
        RECT 4.400 1238.600 1496.000 1240.000 ;
        RECT 4.000 880.960 1496.000 1238.600 ;
        RECT 4.000 879.560 1495.600 880.960 ;
        RECT 4.000 619.840 1496.000 879.560 ;
        RECT 4.400 618.440 1496.000 619.840 ;
        RECT 4.000 260.800 1496.000 618.440 ;
        RECT 4.000 259.400 1495.600 260.800 ;
        RECT 4.000 10.715 1496.000 259.400 ;
      LAYER met4 ;
        RECT 714.240 578.175 788.640 1056.545 ;
        RECT 791.040 578.175 865.440 1056.545 ;
        RECT 867.840 578.175 919.705 1056.545 ;
  END
END user_proj_example
END LIBRARY

