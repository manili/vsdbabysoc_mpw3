VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avsdpll
  CLASS BLOCK ;
  FOREIGN avsdpll ;
  ORIGIN 0.000 0.000 ;
  SIZE 164.380 BY 261.220 ;
  PIN REF
    PORT
      LAYER met2 ;
        RECT 0.010 146.480 58.375 147.670 ;
    END
  END REF
  PIN ENb_VCO
    PORT
      LAYER met2 ;
        RECT 0.010 139.580 112.380 140.920 ;
    END
  END ENb_VCO
  PIN ENb_CP
    PORT
      LAYER met2 ;
        RECT 0.010 135.030 110.000 136.440 ;
    END
  END ENb_CP
  PIN VCO_IN
    PORT
      LAYER met2 ;
        RECT 0.010 105.420 128.280 106.320 ;
    END
  END VCO_IN
  PIN CLK
    PORT
      LAYER met2 ;
        RECT 0.010 108.550 119.280 110.220 ;
    END
  END CLK
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 159.950 3.655 164.380 257.605 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.220 14.855 150.650 245.265 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 50.130 113.170 125.650 144.880 ;
      LAYER met1 ;
        RECT 0.010 113.170 125.720 145.400 ;
      LAYER met2 ;
        RECT 58.655 146.200 128.280 147.690 ;
        RECT 0.070 141.200 128.280 146.200 ;
        RECT 112.660 139.300 128.280 141.200 ;
        RECT 0.070 136.720 128.280 139.300 ;
        RECT 110.280 134.750 128.280 136.720 ;
        RECT 0.070 110.500 128.280 134.750 ;
        RECT 119.560 108.270 128.280 110.500 ;
        RECT 0.070 106.600 128.280 108.270 ;
      LAYER met3 ;
        RECT 0.000 0.000 164.380 261.220 ;
      LAYER met4 ;
        RECT 0.010 258.005 164.380 261.220 ;
        RECT 0.010 245.665 159.550 258.005 ;
        RECT 0.010 14.455 145.820 245.665 ;
        RECT 151.050 14.455 159.550 245.665 ;
        RECT 0.010 3.255 159.550 14.455 ;
        RECT 0.010 0.000 164.380 3.255 ;
  END
END avsdpll
END LIBRARY

