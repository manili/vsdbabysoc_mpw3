VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avsddac
  CLASS BLOCK ;
  FOREIGN avsddac ;
  ORIGIN 0.000 0.000 ;
  SIZE 1520.000 BY 1110.070 ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.150 1109.500 169.650 1110.000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.450 1109.500 184.950 1110.000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.000 1109.500 202.500 1110.000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.610 1109.500 456.110 1110.000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.340 1109.500 233.840 1110.000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.380 1109.500 351.880 1110.000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.700 0.000 1034.200 0.500 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.070 0.000 1089.570 0.500 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.460 0.000 1140.960 0.500 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.950 0.000 1174.450 0.500 ;
    END
  END D[9]
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.150 1109.500 1187.650 1110.000 ;
    END
  END OUT
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1410.000 229.110 1460.000 880.790 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1470.000 169.070 1520.000 940.740 ;
    END
  END vccd1
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.120 1109.570 166.620 1110.070 ;
    END
  END VREFH
  PIN VREFL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.940 60.000 990.440 60.500 ;
    END
  END VREFL
  OBS
      LAYER li1 ;
        RECT 160.000 280.000 1187.420 1110.000 ;
      LAYER met1 ;
        RECT 163.980 0.000 1336.590 1110.070 ;
      LAYER met2 ;
        RECT 60.000 308.860 1188.610 839.130 ;
      LAYER met3 ;
        RECT 0.000 120.000 1520.000 990.000 ;
      LAYER met4 ;
        RECT 0.000 941.140 1520.000 990.000 ;
        RECT 0.000 881.190 1469.600 941.140 ;
        RECT 0.000 228.710 1409.600 881.190 ;
        RECT 1460.400 228.710 1469.600 881.190 ;
        RECT 0.000 168.670 1469.600 228.710 ;
        RECT 0.000 120.000 1520.000 168.670 ;
  END
END avsddac
END LIBRARY

